library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity nco8 is
	port (
		i_clk			: in std_logic;
		i_clk_rst		: in std_logic;
		i_fcw			: in std_logic_vector(7 downto 0);
		o_nco			: out std_logic_vector(7 downto 0)
	);
end entity;

architecture RTL of nco8 is 

	type sine_LUT_type is array (0 to 255) of std_logic_vector (7 downto 0);
	
	constant sine_lut : sine_LUT_type := (
		"10000000", -- LUT[0] == 128
		"10000011", -- LUT[1] == 131
		"10000110", -- LUT[2] == 134
		"10001001", -- LUT[3] == 137
		"10001100", -- LUT[4] == 140
		"10001111", -- LUT[5] == 143
		"10010010", -- LUT[6] == 146
		"10010101", -- LUT[7] == 149
		"10011000", -- LUT[8] == 152
		"10011011", -- LUT[9] == 155
		"10011110", -- LUT[10] == 158
		"10100010", -- LUT[11] == 162
		"10100101", -- LUT[12] == 165
		"10100111", -- LUT[13] == 167
		"10101010", -- LUT[14] == 170
		"10101101", -- LUT[15] == 173
		"10110000", -- LUT[16] == 176
		"10110011", -- LUT[17] == 179
		"10110110", -- LUT[18] == 182
		"10111001", -- LUT[19] == 185
		"10111100", -- LUT[20] == 188
		"10111110", -- LUT[21] == 190
		"11000001", -- LUT[22] == 193
		"11000100", -- LUT[23] == 196
		"11000110", -- LUT[24] == 198
		"11001001", -- LUT[25] == 201
		"11001011", -- LUT[26] == 203
		"11001110", -- LUT[27] == 206
		"11010000", -- LUT[28] == 208
		"11010011", -- LUT[29] == 211
		"11010101", -- LUT[30] == 213
		"11010111", -- LUT[31] == 215
		"11011010", -- LUT[32] == 218
		"11011100", -- LUT[33] == 220
		"11011110", -- LUT[34] == 222
		"11100000", -- LUT[35] == 224
		"11100010", -- LUT[36] == 226
		"11100100", -- LUT[37] == 228
		"11100110", -- LUT[38] == 230
		"11101000", -- LUT[39] == 232
		"11101010", -- LUT[40] == 234
		"11101011", -- LUT[41] == 235
		"11101101", -- LUT[42] == 237
		"11101110", -- LUT[43] == 238
		"11110000", -- LUT[44] == 240
		"11110001", -- LUT[45] == 241
		"11110011", -- LUT[46] == 243
		"11110100", -- LUT[47] == 244
		"11110101", -- LUT[48] == 245
		"11110110", -- LUT[49] == 246
		"11111000", -- LUT[50] == 248
		"11111001", -- LUT[51] == 249
		"11111010", -- LUT[52] == 250
		"11111010", -- LUT[53] == 250
		"11111011", -- LUT[54] == 251
		"11111100", -- LUT[55] == 252
		"11111101", -- LUT[56] == 253
		"11111101", -- LUT[57] == 253
		"11111110", -- LUT[58] == 254
		"11111110", -- LUT[59] == 254
		"11111110", -- LUT[60] == 254
		"11111111", -- LUT[61] == 255
		"11111111", -- LUT[62] == 255
		"11111111", -- LUT[63] == 255
		"11111111", -- LUT[64] == 255
		"11111111", -- LUT[65] == 255
		"11111111", -- LUT[66] == 255
		"11111111", -- LUT[67] == 255
		"11111110", -- LUT[68] == 254
		"11111110", -- LUT[69] == 254
		"11111110", -- LUT[70] == 254
		"11111101", -- LUT[71] == 253
		"11111101", -- LUT[72] == 253
		"11111100", -- LUT[73] == 252
		"11111011", -- LUT[74] == 251
		"11111010", -- LUT[75] == 250
		"11111010", -- LUT[76] == 250
		"11111001", -- LUT[77] == 249
		"11111000", -- LUT[78] == 248
		"11110110", -- LUT[79] == 246
		"11110101", -- LUT[80] == 245
		"11110100", -- LUT[81] == 244
		"11110011", -- LUT[82] == 243
		"11110001", -- LUT[83] == 241
		"11110000", -- LUT[84] == 240
		"11101110", -- LUT[85] == 238
		"11101101", -- LUT[86] == 237
		"11101011", -- LUT[87] == 235
		"11101010", -- LUT[88] == 234
		"11101000", -- LUT[89] == 232
		"11100110", -- LUT[90] == 230
		"11100100", -- LUT[91] == 228
		"11100010", -- LUT[92] == 226
		"11100000", -- LUT[93] == 224
		"11011110", -- LUT[94] == 222
		"11011100", -- LUT[95] == 220
		"11011010", -- LUT[96] == 218
		"11010111", -- LUT[97] == 215
		"11010101", -- LUT[98] == 213
		"11010011", -- LUT[99] == 211
		"11010000", -- LUT[100] == 208
		"11001110", -- LUT[101] == 206
		"11001011", -- LUT[102] == 203
		"11001001", -- LUT[103] == 201
		"11000110", -- LUT[104] == 198
		"11000100", -- LUT[105] == 196
		"11000001", -- LUT[106] == 193
		"10111110", -- LUT[107] == 190
		"10111100", -- LUT[108] == 188
		"10111001", -- LUT[109] == 185
		"10110110", -- LUT[110] == 182
		"10110011", -- LUT[111] == 179
		"10110000", -- LUT[112] == 176
		"10101101", -- LUT[113] == 173
		"10101010", -- LUT[114] == 170
		"10100111", -- LUT[115] == 167
		"10100101", -- LUT[116] == 165
		"10100010", -- LUT[117] == 162
		"10011110", -- LUT[118] == 158
		"10011011", -- LUT[119] == 155
		"10011000", -- LUT[120] == 152
		"10010101", -- LUT[121] == 149
		"10010010", -- LUT[122] == 146
		"10001111", -- LUT[123] == 143
		"10001100", -- LUT[124] == 140
		"10001001", -- LUT[125] == 137
		"10000110", -- LUT[126] == 134
		"10000011", -- LUT[127] == 131
		"10000000", -- LUT[128] == 128
		"01111100", -- LUT[129] == 124
		"01111001", -- LUT[130] == 121
		"01110110", -- LUT[131] == 118
		"01110011", -- LUT[132] == 115
		"01110000", -- LUT[133] == 112
		"01101101", -- LUT[134] == 109
		"01101010", -- LUT[135] == 106
		"01100111", -- LUT[136] == 103
		"01100100", -- LUT[137] == 100
		"01100001", -- LUT[138] == 97
		"01011101", -- LUT[139] == 93
		"01011010", -- LUT[140] == 90
		"01011000", -- LUT[141] == 88
		"01010101", -- LUT[142] == 85
		"01010010", -- LUT[143] == 82
		"01001111", -- LUT[144] == 79
		"01001100", -- LUT[145] == 76
		"01001001", -- LUT[146] == 73
		"01000110", -- LUT[147] == 70
		"01000011", -- LUT[148] == 67
		"01000001", -- LUT[149] == 65
		"00111110", -- LUT[150] == 62
		"00111011", -- LUT[151] == 59
		"00111001", -- LUT[152] == 57
		"00110110", -- LUT[153] == 54
		"00110100", -- LUT[154] == 52
		"00110001", -- LUT[155] == 49
		"00101111", -- LUT[156] == 47
		"00101100", -- LUT[157] == 44
		"00101010", -- LUT[158] == 42
		"00101000", -- LUT[159] == 40
		"00100101", -- LUT[160] == 37
		"00100011", -- LUT[161] == 35
		"00100001", -- LUT[162] == 33
		"00011111", -- LUT[163] == 31
		"00011101", -- LUT[164] == 29
		"00011011", -- LUT[165] == 27
		"00011001", -- LUT[166] == 25
		"00010111", -- LUT[167] == 23
		"00010101", -- LUT[168] == 21
		"00010100", -- LUT[169] == 20
		"00010010", -- LUT[170] == 18
		"00010001", -- LUT[171] == 17
		"00001111", -- LUT[172] == 15
		"00001110", -- LUT[173] == 14
		"00001100", -- LUT[174] == 12
		"00001011", -- LUT[175] == 11
		"00001010", -- LUT[176] == 10
		"00001001", -- LUT[177] == 9
		"00000111", -- LUT[178] == 7
		"00000110", -- LUT[179] == 6
		"00000101", -- LUT[180] == 5
		"00000101", -- LUT[181] == 5
		"00000100", -- LUT[182] == 4
		"00000011", -- LUT[183] == 3
		"00000010", -- LUT[184] == 2
		"00000010", -- LUT[185] == 2
		"00000001", -- LUT[186] == 1
		"00000001", -- LUT[187] == 1
		"00000001", -- LUT[188] == 1
		"00000000", -- LUT[189] == 0
		"00000000", -- LUT[190] == 0
		"00000000", -- LUT[191] == 0
		"00000000", -- LUT[192] == 0
		"00000000", -- LUT[193] == 0
		"00000000", -- LUT[194] == 0
		"00000000", -- LUT[195] == 0
		"00000001", -- LUT[196] == 1
		"00000001", -- LUT[197] == 1
		"00000001", -- LUT[198] == 1
		"00000010", -- LUT[199] == 2
		"00000010", -- LUT[200] == 2
		"00000011", -- LUT[201] == 3
		"00000100", -- LUT[202] == 4
		"00000101", -- LUT[203] == 5
		"00000101", -- LUT[204] == 5
		"00000110", -- LUT[205] == 6
		"00000111", -- LUT[206] == 7
		"00001001", -- LUT[207] == 9
		"00001010", -- LUT[208] == 10
		"00001011", -- LUT[209] == 11
		"00001100", -- LUT[210] == 12
		"00001110", -- LUT[211] == 14
		"00001111", -- LUT[212] == 15
		"00010001", -- LUT[213] == 17
		"00010010", -- LUT[214] == 18
		"00010100", -- LUT[215] == 20
		"00010101", -- LUT[216] == 21
		"00010111", -- LUT[217] == 23
		"00011001", -- LUT[218] == 25
		"00011011", -- LUT[219] == 27
		"00011101", -- LUT[220] == 29
		"00011111", -- LUT[221] == 31
		"00100001", -- LUT[222] == 33
		"00100011", -- LUT[223] == 35
		"00100101", -- LUT[224] == 37
		"00101000", -- LUT[225] == 40
		"00101010", -- LUT[226] == 42
		"00101100", -- LUT[227] == 44
		"00101111", -- LUT[228] == 47
		"00110001", -- LUT[229] == 49
		"00110100", -- LUT[230] == 52
		"00110110", -- LUT[231] == 54
		"00111001", -- LUT[232] == 57
		"00111011", -- LUT[233] == 59
		"00111110", -- LUT[234] == 62
		"01000001", -- LUT[235] == 65
		"01000011", -- LUT[236] == 67
		"01000110", -- LUT[237] == 70
		"01001001", -- LUT[238] == 73
		"01001100", -- LUT[239] == 76
		"01001111", -- LUT[240] == 79
		"01010010", -- LUT[241] == 82
		"01010101", -- LUT[242] == 85
		"01011000", -- LUT[243] == 88
		"01011010", -- LUT[244] == 90
		"01011101", -- LUT[245] == 93
		"01100001", -- LUT[246] == 97
		"01100100", -- LUT[247] == 100
		"01100111", -- LUT[248] == 103
		"01101010", -- LUT[249] == 106
		"01101101", -- LUT[250] == 109
		"01110000", -- LUT[251] == 112
		"01110011", -- LUT[252] == 115
		"01110110", -- LUT[253] == 118
		"01111001", -- LUT[254] == 121
		"01111100"  -- LUT[255] == 124
	);

	signal r_phase 		: unsigned(7 downto 0) := (others => '0');

	begin
		process (i_clk, i_clk_rst)
    	begin
			
			if(rising_edge(i_clk)) then
				if(i_clk_rst = '1') then
					r_phase <= (others => '0');
				end if;
				r_phase <= r_phase + unsigned(i_fcw);
				o_nco <= sine_lut(to_integer(r_phase));
			end if;
		end process;
		
end RTL;
		